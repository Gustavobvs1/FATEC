<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>17.2411,44.248,223.527,-58.4509</PageViewport>
<gate>
<ID>4</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>148,-0.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>6 </input>
<input>
<ID>IN_4</ID>4 </input>
<input>
<ID>IN_5</ID>3 </input>
<input>
<ID>IN_6</ID>2 </input>
<input>
<ID>IN_7</ID>1 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_DFF_LOW</type>
<position>111,-20</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>6 </output>
<input>
<ID>clock</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_DFF_LOW</type>
<position>111,-29.5</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>7 </output>
<input>
<ID>clock</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_DFF_LOW</type>
<position>111,-41</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>8 </output>
<input>
<ID>clock</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_DFF_LOW</type>
<position>111.5,-52</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>9 </output>
<input>
<ID>clock</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>102,-18</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>102,-27</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>100.5,-38.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>101,-49.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>58</ID>
<type>AE_DFF_LOW</type>
<position>111,-11</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>4 </output>
<input>
<ID>clock</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_DFF_LOW</type>
<position>113,-2.5</position>
<input>
<ID>IN_0</ID>25 </input>
<output>
<ID>OUT_0</ID>3 </output>
<input>
<ID>clock</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_DFF_LOW</type>
<position>111.5,6.5</position>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>2 </output>
<input>
<ID>clock</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_DFF_LOW</type>
<position>115,16</position>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>1 </output>
<input>
<ID>clock</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>105,18</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_TOGGLE</type>
<position>103.5,8.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>65.5,-11</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>103.5,-1</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>103,-8.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118,18,143,18</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>143 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>143,3.5,143,18</points>
<connection>
<GID>4</GID>
<name>IN_7</name></connection>
<intersection>18 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,2.5,128.5,9</points>
<intersection>2.5 1</intersection>
<intersection>9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,2.5,143,2.5</points>
<connection>
<GID>4</GID>
<name>IN_6</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,9,128.5,9</points>
<intersection>114.5 3</intersection>
<intersection>128.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114.5,8.5,114.5,9</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>9 2</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-0.5,129.5,1.5</points>
<intersection>-0.5 2</intersection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,1.5,143,1.5</points>
<connection>
<GID>4</GID>
<name>IN_5</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-0.5,129.5,-0.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-9,134,0.5</points>
<intersection>-9 2</intersection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,0.5,143,0.5</points>
<connection>
<GID>4</GID>
<name>IN_4</name></connection>
<intersection>134 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-9,134,-9</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>134 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-18,135,-0.5</points>
<intersection>-18 2</intersection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-0.5,143,-0.5</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-18,135,-18</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-27.5,136,-1.5</points>
<intersection>-27.5 2</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-1.5,143,-1.5</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-27.5,136,-27.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-39,137,-2.5</points>
<intersection>-39 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137,-2.5,143,-2.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-39,137,-39</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-50,138,-3.5</points>
<intersection>-50 2</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-3.5,143,-3.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-50,138,-50</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-18,108,-18</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-39,105,-38.5</points>
<intersection>-39 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-39,108,-39</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102.5,-38.5,105,-38.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-50,105.5,-49.5</points>
<intersection>-50 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-50,108.5,-50</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-49.5,105.5,-49.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-27.5,106,-27</points>
<intersection>-27.5 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-27.5,108,-27.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-27,106,-27</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-11,77,15</points>
<intersection>-11 2</intersection>
<intersection>15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,15,112,15</points>
<connection>
<GID>64</GID>
<name>clock</name></connection>
<intersection>77 0</intersection>
<intersection>90.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>67.5,-11,77,-11</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>77 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>90.5,-53,90.5,15</points>
<intersection>-53 16</intersection>
<intersection>-42 14</intersection>
<intersection>-30.5 12</intersection>
<intersection>-21 10</intersection>
<intersection>-12 8</intersection>
<intersection>-3.5 6</intersection>
<intersection>5.5 4</intersection>
<intersection>15 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>90.5,5.5,108.5,5.5</points>
<connection>
<GID>62</GID>
<name>clock</name></connection>
<intersection>90.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>90.5,-3.5,110,-3.5</points>
<connection>
<GID>60</GID>
<name>clock</name></connection>
<intersection>90.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>90.5,-12,108,-12</points>
<connection>
<GID>58</GID>
<name>clock</name></connection>
<intersection>90.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>90.5,-21,108,-21</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<intersection>90.5 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>90.5,-30.5,108,-30.5</points>
<connection>
<GID>8</GID>
<name>clock</name></connection>
<intersection>90.5 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>90.5,-42,108,-42</points>
<connection>
<GID>10</GID>
<name>clock</name></connection>
<intersection>90.5 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>90.5,-53,108.5,-53</points>
<connection>
<GID>12</GID>
<name>clock</name></connection>
<intersection>90.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107,18,112,18</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105.5,8.5,108.5,8.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-1,107.5,-0.5</points>
<intersection>-1 2</intersection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-0.5,110,-0.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,-1,107.5,-1</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-8.5,108,-8.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>108 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>108,-9,108,-8.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-0.000499424,322.623,1394,-371.377</PageViewport></page 1>
<page 2>
<PageViewport>-0.000499424,322.623,1394,-371.377</PageViewport></page 2>
<page 3>
<PageViewport>-0.000499424,322.623,1394,-371.377</PageViewport></page 3>
<page 4>
<PageViewport>-0.000499424,322.623,1394,-371.377</PageViewport></page 4>
<page 5>
<PageViewport>-0.000499424,322.623,1394,-371.377</PageViewport></page 5>
<page 6>
<PageViewport>-0.000499424,322.623,1394,-371.377</PageViewport></page 6>
<page 7>
<PageViewport>-0.000499424,322.623,1394,-371.377</PageViewport></page 7>
<page 8>
<PageViewport>-0.000499424,322.623,1394,-371.377</PageViewport></page 8>
<page 9>
<PageViewport>-0.000499424,322.623,1394,-371.377</PageViewport></page 9></circuit>