<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-978.507,582.34,-765.337,476.214</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>2.5,-14</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>-903.5,503</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>9.5,-13.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>-901.5,497</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-878,509.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>7 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>-817.5,507.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>-812,502.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>41,-22</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>-889.5,561</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_AND2</type>
<position>-889.5,554.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>3,-18</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND2</type>
<position>-889.5,547</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>10,-18</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND3</type>
<position>-877.5,554.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<input>
<ID>IN_2</ID>5 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>20</ID>
<type>AI_XOR2</type>
<position>-889.5,571.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AI_XOR2</type>
<position>-876,567.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-849,567.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<input>
<ID>IN_2</ID>33 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND2</type>
<position>-839,540</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AI_XOR2</type>
<position>-854,545.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-821.5,522</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>11 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>26</ID>
<type>AI_XOR2</type>
<position>29,-21</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>AI_XOR2</type>
<position>38.5,-26</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_AND2</type>
<position>30,-31.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_AND2</type>
<position>30,-38.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_AND2</type>
<position>30,-44.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>AE_OR3</type>
<position>43,-37.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>19 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>19,-18</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>19.5,-13.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>49,-26</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>GA_LED</type>
<position>51,-37.5</position>
<input>
<ID>N_in0</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>24,40</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_TOGGLE</type>
<position>26.5,35.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>28,31.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>71</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>51.5,39</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>72</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>97.5,45</position>
<input>
<ID>IN_3</ID>2 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>74</ID>
<type>AI_XOR2</type>
<position>34,65.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AI_XOR2</type>
<position>42.5,61.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>61.5,66.5</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_AND2</type>
<position>34.5,55.5</position>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_AND2</type>
<position>34.5,50</position>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_AND2</type>
<position>34.5,45</position>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AE_OR3</type>
<position>44.5,50</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>38 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_OR2</type>
<position>66,52.5</position>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_AND2</type>
<position>74.5,47</position>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>88</ID>
<type>AI_XOR2</type>
<position>87,73.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>AI_XOR2</type>
<position>99,68.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_AND2</type>
<position>99.5,63</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_AND2</type>
<position>100,58</position>
<input>
<ID>IN_1</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AA_AND2</type>
<position>100.5,53</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_TOGGLE</type>
<position>105,39.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_TOGGLE</type>
<position>107,34.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_TOGGLE</type>
<position>109,29</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,31.5,87,54</points>
<intersection>31.5 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,31.5,87,31.5</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87,54,97.5,54</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,29,89,52</points>
<intersection>29 1</intersection>
<intersection>47 3</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89,29,107,29</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,52,97.5,52</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>89 0</intersection>
<intersection>92.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>89,47,94.5,47</points>
<connection>
<GID>72</GID>
<name>IN_3</name></connection>
<intersection>89 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>92.5,52,92.5,69.5</points>
<intersection>52 2</intersection>
<intersection>69.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>92.5,69.5,96,69.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>92.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-883.5,556.5,-883.5,561</points>
<intersection>556.5 1</intersection>
<intersection>561 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-883.5,556.5,-880.5,556.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-883.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-886.5,561,-883.5,561</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>-883.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-886.5,554.5,-880.5,554.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>-886.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-886.5,554.5,-886.5,554.5</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>554.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-883.5,547,-883.5,552.5</points>
<intersection>547 2</intersection>
<intersection>552.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-883.5,552.5,-880.5,552.5</points>
<connection>
<GID>18</GID>
<name>IN_2</name></connection>
<intersection>-883.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-886.5,547,-883.5,547</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>-883.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-900,503,-900,570.5</points>
<intersection>503 1</intersection>
<intersection>509.5 6</intersection>
<intersection>548 4</intersection>
<intersection>562 5</intersection>
<intersection>570.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-901.5,503,-900,503</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-900 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-900,570.5,-892.5,570.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-900 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-900,548,-892.5,548</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-900 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-900,562,-892.5,562</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-900 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-900,509.5,-881,509.5</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>-900 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-906,502.5,-906,572.5</points>
<intersection>502.5 2</intersection>
<intersection>546 8</intersection>
<intersection>555.5 3</intersection>
<intersection>572.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-906,572.5,-892.5,572.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-906 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-906,502.5,-814,502.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>-906 0</intersection>
<intersection>-830.5 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-906,555.5,-892.5,555.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-906 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-830.5,502.5,-830.5,522</points>
<intersection>502.5 2</intersection>
<intersection>522 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-830.5,522,-824.5,522</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>-830.5 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-906,546,-892.5,546</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>-906 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-25,33.5,-21</points>
<intersection>-25 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-25,35.5,-25</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-21,33.5,-21</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-897.5,551,-897.5,566.5</points>
<intersection>551 2</intersection>
<intersection>553.5 4</intersection>
<intersection>560 3</intersection>
<intersection>566.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-897.5,566.5,-879,566.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>-897.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-897.5,551,-839,551</points>
<intersection>-897.5 0</intersection>
<intersection>-839 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-897.5,560,-892.5,560</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>-897.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-897.5,553.5,-892.5,553.5</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>-897.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-839,543,-839,551</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<intersection>551 2</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-882.5,568.5,-882.5,571.5</points>
<intersection>568.5 1</intersection>
<intersection>571.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-882.5,568.5,-879,568.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-882.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-886.5,571.5,-882.5,571.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>-882.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-35.5,36.5,-31.5</points>
<intersection>-35.5 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-35.5,40,-35.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-31.5,36.5,-31.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-38.5,36.5,-37.5</points>
<intersection>-38.5 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-37.5,40,-37.5</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-38.5,36.5,-38.5</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-44.5,36.5,-39.5</points>
<intersection>-44.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-39.5,40,-39.5</points>
<connection>
<GID>39</GID>
<name>IN_2</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-44.5,36.5,-44.5</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-45.5,5,-18</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-45.5 1</intersection>
<intersection>-37.5 3</intersection>
<intersection>-20 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-45.5,27,-45.5</points>
<connection>
<GID>33</GID>
<name>IN_1</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>5,-37.5,27,-37.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>5,-20,26,-20</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-43.5,14,-18</points>
<intersection>-43.5 1</intersection>
<intersection>-30.5 3</intersection>
<intersection>-22 5</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-43.5,27,-43.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-18,14,-18</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>14,-30.5,27,-30.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>14,-22,26,-22</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-39.5,24,-18</points>
<intersection>-39.5 1</intersection>
<intersection>-32.5 3</intersection>
<intersection>-27 5</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-39.5,27,-39.5</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-18,24,-18</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24,-32.5,27,-32.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>24,-27,35.5,-27</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41.5,-26,48,-26</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,-37.5,50,-37.5</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<connection>
<GID>47</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-851,497,-851,542.5</points>
<intersection>497 1</intersection>
<intersection>529.5 3</intersection>
<intersection>542.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-899.5,497,-851,497</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>-881 6</intersection>
<intersection>-851 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-853,542.5,-851,542.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>-851 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-851,529.5,-838,529.5</points>
<intersection>-851 0</intersection>
<intersection>-838 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-838,529.5,-838,537</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>529.5 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-881,497,-881,508.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>497 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-855,507.5,-855,542.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>507.5 1</intersection>
<intersection>531.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-855,507.5,-819.5,507.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-855 0</intersection>
<intersection>-825 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-825,507.5,-825,521</points>
<intersection>507.5 1</intersection>
<intersection>521 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-855,531.5,-840,531.5</points>
<intersection>-855 0</intersection>
<intersection>-840 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-840,531.5,-840,537</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>531.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-825,521,-824.5,521</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-825 2</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-852,548.5,-852,566.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>548.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-854,548.5,-852,548.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>-852 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-873,567.5,-852,567.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<connection>
<GID>21</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-863,554.5,-863,568.5</points>
<intersection>554.5 2</intersection>
<intersection>568.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-863,568.5,-852,568.5</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>-863 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-874.5,554.5,-863,554.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>-863 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,52,39.5,55.5</points>
<intersection>52 1</intersection>
<intersection>55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,52,41.5,52</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,55.5,39.5,55.5</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,50,41.5,50</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<connection>
<GID>79</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,45,39.5,48</points>
<intersection>45 2</intersection>
<intersection>48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,48,41.5,48</points>
<connection>
<GID>82</GID>
<name>IN_2</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,45,39.5,45</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,50,87,67.5</points>
<intersection>50 2</intersection>
<intersection>57 3</intersection>
<intersection>67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,67.5,96,67.5</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47.5,50,87,50</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>87,57,97,57</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,33.4057,384.138,-157.837</PageViewport></page 1>
<page 2>
<PageViewport>0,33.4057,384.138,-157.837</PageViewport></page 2>
<page 3>
<PageViewport>0,33.4057,384.138,-157.837</PageViewport></page 3>
<page 4>
<PageViewport>0,33.4057,384.138,-157.837</PageViewport></page 4>
<page 5>
<PageViewport>0,33.4057,384.138,-157.837</PageViewport></page 5>
<page 6>
<PageViewport>0,33.4057,384.138,-157.837</PageViewport></page 6>
<page 7>
<PageViewport>0,33.4057,384.138,-157.837</PageViewport></page 7>
<page 8>
<PageViewport>0,33.4057,384.138,-157.837</PageViewport></page 8>
<page 9>
<PageViewport>0,33.4057,384.138,-157.837</PageViewport></page 9></circuit>