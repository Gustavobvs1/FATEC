<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-878.068,584.842,-665.347,478.939</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>-823.5,563.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-825,533.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>-712.5,537.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>BE_JKFF_LOW</type>
<position>-789,551.5</position>
<input>
<ID>J</ID>3 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>5 </output>
<input>
<ID>clock</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>BE_JKFF_LOW</type>
<position>-753,546.5</position>
<input>
<ID>J</ID>7 </input>
<input>
<ID>K</ID>6 </input>
<output>
<ID>Q</ID>8 </output>
<input>
<ID>clock</ID>12 </input>
<output>
<ID>nQ</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_OR2</type>
<position>-805.5,552</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_SMALL_INVERTER</type>
<position>-810.5,553</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>-716.5,537.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>-769,552</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_SMALL_INVERTER</type>
<position>-759,545</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-797,549.5,-797,552</points>
<intersection>549.5 1</intersection>
<intersection>552 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-797,549.5,-792,549.5</points>
<connection>
<GID>8</GID>
<name>K</name></connection>
<intersection>-797 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-802.5,552,-797,552</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>-797 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-821.5,563.5,-776,563.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-812.5 3</intersection>
<intersection>-792 5</intersection>
<intersection>-776 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-812.5,553,-812.5,563.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>563.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-776,545,-776,563.5</points>
<intersection>545 6</intersection>
<intersection>553 7</intersection>
<intersection>563.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-792,553.5,-792,563.5</points>
<connection>
<GID>8</GID>
<name>J</name></connection>
<intersection>563.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-776,545,-761,545</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-776 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-776,553,-772,553</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-776 4</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-808.5,553,-808.5,553</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-779,551,-779,553.5</points>
<intersection>551 1</intersection>
<intersection>553.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-779,551,-772,551</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>-779 0</intersection>
<intersection>-778.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-786,553.5,-779,553.5</points>
<connection>
<GID>8</GID>
<name>Q</name></connection>
<intersection>-779 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-778.5,536.5,-778.5,551</points>
<intersection>536.5 4</intersection>
<intersection>551 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-778.5,536.5,-719.5,536.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>-778.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-757,544.5,-757,545</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>544.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-757,544.5,-756,544.5</points>
<connection>
<GID>10</GID>
<name>K</name></connection>
<intersection>-757 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-761,548.5,-761,552</points>
<intersection>548.5 1</intersection>
<intersection>552 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-761,548.5,-756,548.5</points>
<connection>
<GID>10</GID>
<name>J</name></connection>
<intersection>-761 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-766,552,-761,552</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>-761 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-734.5,538.5,-734.5,548.5</points>
<intersection>538.5 1</intersection>
<intersection>548.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-734.5,538.5,-719.5,538.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-734.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-750,548.5,-734.5,548.5</points>
<connection>
<GID>10</GID>
<name>Q</name></connection>
<intersection>-734.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-713.5,537.5,-713.5,537.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>6</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-808.5,540.5,-750,540.5</points>
<intersection>-808.5 4</intersection>
<intersection>-750 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-750,540.5,-750,544.5</points>
<connection>
<GID>10</GID>
<name>nQ</name></connection>
<intersection>540.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-808.5,540.5,-808.5,551</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>540.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-823,533.5,-756,533.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-792 4</intersection>
<intersection>-756 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-756,533.5,-756,546.5</points>
<connection>
<GID>10</GID>
<name>clock</name></connection>
<intersection>533.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-792,533.5,-792,551.5</points>
<connection>
<GID>8</GID>
<name>clock</name></connection>
<intersection>533.5 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,138.544,1211.51,-464.605</PageViewport></page 1>
<page 2>
<PageViewport>0,138.544,1211.51,-464.605</PageViewport></page 2>
<page 3>
<PageViewport>0,138.544,1211.51,-464.605</PageViewport></page 3>
<page 4>
<PageViewport>0,138.544,1211.51,-464.605</PageViewport></page 4>
<page 5>
<PageViewport>0,138.544,1211.51,-464.605</PageViewport></page 5>
<page 6>
<PageViewport>0,138.544,1211.51,-464.605</PageViewport></page 6>
<page 7>
<PageViewport>0,138.544,1211.51,-464.605</PageViewport></page 7>
<page 8>
<PageViewport>0,138.544,1211.51,-464.605</PageViewport></page 8>
<page 9>
<PageViewport>0,138.544,1211.51,-464.605</PageViewport></page 9></circuit>